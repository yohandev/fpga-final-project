`default_nettype none

module top_level(
    input wire clk_100mhz,
    
    input wire [15:0]   sw,
    input wire [3:0]    btn
);

// wow, so empty

endmodule

`default_nettype wire