`ifndef FIXED_SV
`define FIXED_SV

typedef struct packed {
    logic signed [31:0] inner;
} fixed;

// Number of bits in the decimal portion of fixed numbers
parameter D = 15;

`define fadd(a, b) fixed'(signed'(a) + signed'(b))
`define fsub(a, b) fixed'(signed'(a) - signed'(b))
`define fmul(a, b) fixed'(32'((64'(signed'(a)) * 64'(signed'(b))) >>> D))

`define FIXED_1 fixed'(32'sh8000)
`define FIXED_1_5 fixed'(32'shC000)

module fixed_inv_sqrt(
    input wire clk_in,

    input fixed in,
    output fixed out
);
    fixed lut;

    always_comb begin
        // Generated with fixed_inv_sqrt.py [D=15]
        unique casez (in)
            32'sb?01?????????????????????????????: lut = 32'sh93;
            32'sb?001????????????????????????????: lut = 32'shd1;
            32'sb?0001???????????????????????????: lut = 32'sh127;
            32'sb?00001??????????????????????????: lut = 32'sh1a2;
            32'sb?000001?????????????????????????: lut = 32'sh24f;
            32'sb?0000001????????????????????????: lut = 32'sh344;
            32'sb?00000001???????????????????????: lut = 32'sh49e;
            32'sb?000000001??????????????????????: lut = 32'sh688;
            32'sb?0000000001?????????????????????: lut = 32'sh93c;
            32'sb?00000000001????????????????????: lut = 32'shd10;
            32'sb?000000000001???????????????????: lut = 32'sh1279;
            32'sb?0000000000001??????????????????: lut = 32'sh1a20;
            32'sb?00000000000001?????????????????: lut = 32'sh24f3;
            32'sb?000000000000001????????????????: lut = 32'sh3441;
            32'sb?0000000000000001???????????????: lut = 32'sh49e6;
            32'sb?00000000000000001??????????????: lut = 32'sh6882;
            32'sb?000000000000000001?????????????: lut = 32'sh93cd;
            32'sb?0000000000000000001????????????: lut = 32'shd105;
            32'sb?00000000000000000001???????????: lut = 32'sh1279a;
            32'sb?000000000000000000001??????????: lut = 32'sh1a20b;
            32'sb?0000000000000000000001?????????: lut = 32'sh24f34;
            32'sb?00000000000000000000001????????: lut = 32'sh34417;
            32'sb?000000000000000000000001???????: lut = 32'sh49e69;
            32'sb?0000000000000000000000001??????: lut = 32'sh6882f;
            32'sb?00000000000000000000000001?????: lut = 32'sh93cd3;
            32'sb?000000000000000000000000001????: lut = 32'shd105e;
            32'sb?0000000000000000000000000001???: lut = 32'sh1279a7;
            32'sb?00000000000000000000000000001??: lut = 32'sh1a20bd;
            32'sb?000000000000000000000000000001?: lut = 32'sh24f34e;
            32'sb?0000000000000000000000000000001: lut = 32'sh34417a;
            default: lut = 32'sh5a8279;
        endcase
    end

    fixed in_pipe0, in_pipe1;
    fixed iter0, iter0_pipe0, iter0_pipe1;
    fixed iter1, iter1_pipe0, iter1_pipe1;

    assign out = iter1;

    always_ff @(posedge clk_in) begin
        // Look-up table
        iter0 <= lut;
        in_pipe0 <= in;

        // Newton's method, first iteration (first intermediate)
        iter1_pipe0 <= `fmul(iter0, iter0);
        iter0_pipe0 <= iter0;
        in_pipe1 <= in_pipe0;

        // Neton's method, first iteration (second intermediate)
        iter0_pipe1 <= iter0_pipe0;
        iter1_pipe1 <= `fmul(fixed'(in_pipe1 >> 1), iter1_pipe0);

        // Newton's method, second iteration (done)
        iter1 <= `fmul(iter0_pipe1, `fsub(`FIXED_1_5, iter1_pipe1));
    end
endmodule

module fixed_testbench(
    input wire clk_in,

    input fixed a,
    input fixed b,

    output fixed add,
    output fixed sub,
    output fixed mul,
    output fixed expr,
    output fixed inv_sqrt
);
    fixed_inv_sqrt fixed_inv_sqrt(
        .clk_in(clk_in),
        .in(a),
        .out(inv_sqrt)
    );

    always_ff @(posedge clk_in) begin
        add <= `fadd(a, b);
        sub <= `fsub(a, b);
        mul <= `fmul(a, b);
        expr <= `fmul(`fadd(`fmul(a, b), `fsub(b, a)), `fsub(a, b));
    end
endmodule

`endif